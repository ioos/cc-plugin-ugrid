netcdf UGRID {
dimensions:
	time   = UNLIMITED ;     // (1 currently)
	nnodes = 5 ;	         // number of nodes
	nedges = 9 ;	         // number of edges
	nfaces = 9 ;             // number of nfaces
    maxnumnodesperface = 7 ; // used for optional connectivities and in fully 3D volume connectivities
	three  = 3 ;             // extraneous dimension, used in face_node_connectivity array
	two    = 2 ;   	         // extraneous dimension, used in edge_node_connectivity array
variables:
  int mesh_topology ;
  	mesh_topology:cf_role                = "mesh_topology" ;
  	mesh_topology:topology_dimension     = 2 ;
  	mesh_topology:edge_dimension         = "nedges" ;
  	mesh_topology:face_dimension         = "nfaces" ;
  	mesh_topology:node_coordinates       = "lon lat" ;
  	mesh_topology:face_coordinates       = "lonc latc" ;
  	mesh_topology:edge_coordinates       = "lone late" ;
    mesh_topology:edge_face_connectivity = "efc" ;
    mesh_topology:edge_node_connectivity = "enc" ;
    mesh_topology:face_edge_connectivity = "fec" ;
  	mesh_topology:face_node_connectivity = "nv" ;
  int mesh_topology2 ;
 	mesh_topology2:cf_role                = "mesh_topology" ;
 	mesh_topology2:topology_dimension     = 2 ;
 	mesh_topology2:edge_dimension         = "nedges" ;
 	mesh_topology2:face_dimension         = "nfaces" ;
 	mesh_topology2:node_coordinates       = "lon lat" ;
 	mesh_topology2:face_coordinates       = "lonc latc" ;
 	mesh_topology2:edge_coordinates       = "lone late" ;
    mesh_topology2:edge_face_connectivity = "efc2" ;
 	mesh_topology2:edge_node_connectivity = "enc2" ;
    mesh_topology2:face_edge_connectivity = "fec2" ;
 	mesh_topology2:face_node_connectivity = "nv2" ;
  int efc(nedges, two) ;                              // edge_face_connectivity array
		efc:long_name   = "edge_face_connectivity" ;
        efc:cf_role     = "edge_face_connectivity" ;
        efc:start_index = 1 ;
        efc:location    = "exists" ;
        efc:mesh        = "mesh_topology" ;
  int efc2(nedges, two) ;                              // edge_face_connectivity array
		efc2:long_name   = "edge_face_connectivity" ;
        efc2:cf_role     = "edge_face_connectivity" ;
        efc2:start_index = 1 ;
        efc2:location    = "exists" ;
        efc2:mesh        = "mesh_topology2" ;
  int enc(nedges, two) ;                              // standard order
		enc:long_name = "edge_node_connectivity" ;
		enc:cf_role = "edge_node_connectivity" ;
		enc:start_index = 1 ;
		enc:location = "exists";
		enc:mesh = "mesh_topology";
  int enc2(nedges, two) ;                              // standard order
		enc2:long_name = "edge_node_connectivity" ;
		enc2:cf_role = "edge_node_connectivity" ;
		enc2:start_index = 1 ;
		enc2:location = "exists";
		enc2:mesh = "mesh_topology2";
  int fec(nfaces, maxnumnodesperface) ;
		fec:long_name    = "face_edge_connectivity" ;
		fec:cf_role      = "face_edge_connectivity" ;
        fec:start_index  = 1 ;
		fec:location     = "exists" ;
		fec:mesh         = "mesh_topology" ;
  int fec2(nfaces, maxnumnodesperface) ;
		fec2:long_name    = "face_edge_connectivity" ;
		fec2:cf_role      = "face_edge_connectivity" ;
        fec2:start_index  = 1 ;
		fec2:location     = "exists" ;
		fec2:mesh         = "mesh_topology2" ;
  float lat(nnodes) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:location = "exists";
		lat:mesh = "mesh_topology";
  float late(nedges) ;
		late:long_name = "latitude centered on edge" ;
		late:standard_name = "latitude" ;
		late:units = "degrees_north" ;
		late:location = "exists";
		late:mesh = "mesh_topology";
  float latc(nfaces) ;
		latc:long_name = "latitude centered on face" ;
		latc:standard_name = "latitude" ;
		latc:units = "degrees_north" ;
		latc:location = "exists";
		latc:mesh = "mesh_topology";
  float lon(nnodes) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:location = "exists";
		lon:mesh = "mesh_topology";
  float lone(nfaces) ;
		lone:long_name = "longitude centered on edge" ;
		lone:standard_name = "longitude" ;
		lone:units = "degrees_east" ;
		lone:location = "exists";
		lone:mesh = "mesh_topology";
  float lonc(nfaces) ;
		lonc:long_name = "longitude centered on face" ;
		lonc:standard_name = "longitude" ;
		lonc:units = "degrees_east" ;
		lonc:location = "exists";
		lonc:mesh = "mesh_topology";
  int nv(three, nfaces) ;                             // nonstandard order
		nv:long_name = "nodes surrounding element" ;
		nv:cf_role = "face_node_connectivity" ;
		nv:start_index = 1 ;
		nv:location = "exists";
		nv:mesh = "mesh_topology";
  int nv2(three, nfaces) ;                            // nonstandard order
		nv2:long_name = "nodes surrounding element" ;
		nv2:cf_role = "face_node_connectivity" ;
		nv2:start_index = 1 ;
		nv2:location = "exists";
		nv2:mesh = "mesh_topology2";
  float temperature(time, nfaces) ;
		temperature:location = "exists";
		temperature:mesh = "mesh_topology";
  float eastward_velocity(time, nnodes) ;
		eastward_velocity:location = "exists";
		eastward_velocity:mesh = "mesh_topology";
  float northward_velocity(time, nnodes) ;
		northward_velocity:location = "exists";
		northward_velocity:mesh = "mesh_topology";
  float flux(time, nedges) ;
		flux:location = "exists" ;
		flux:mesh = "mesh_topology" ;
  int time(time);
		time:standard_name = "time" ;
		time:location = "exists" ;
		time:mesh = "mesh_topology" ;
// global attributes:
		:institution = "School for Marine Science and Technology" ;
		:source = "FVCOM" ;
		:references = "http://fvcom.smast.umassd.edu" ;
		:Conventions = "CF-1.0, UGRID-1.0" ;
}
