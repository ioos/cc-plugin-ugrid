netcdf fvcom_reference {
dimensions:
	time = UNLIMITED ; // (1 currently)
	nele = 8 ;
	node = 4 ;
	siglay = 5 ;
	three = 3 ;
variables:
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1858-11-17 00:00:00" ;
		time:format = "modified julian dat (MJD)" ;
		time:time_zone = "UTC" ;
		time:standard_name = "time" ;
	char Times(time, maxStrlen64) ;
		Times:time_zone = "UTC" ;
	float lon(node) ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(node) ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	float lonc(nele) ;
		lonc:long_name = "Longitude" ;
		lonc:standard_name = "longitude" ;
		lonc:units = "degrees_east" ;
	float latc(nele) ;
		latc:long_name = "Latitude" ;
		latc:standard_name = "latitude" ;
		latc:units = "degrees_north" ;
	float siglay(siglay, node) ;
		siglay:long_name = "Sigma Layers" ;
		siglay:standard_name = "ocean_sigma_coordinate" ;
		siglay:positive = "up" ;
		siglay:valid_min = -1. ;
		siglay:valid_max = 0. ;
		siglay:formula_terms = "sigma: siglay eta: zeta depth: h" ;
	float h(node) ;
		h:long_name = "Bathymetry" ;
		h:standard_name = "sea_floor_depth_below_geoid" ;
		h:units = "m" ;
		h:coordinates = "lat lon" ;
		h:type = "data" ;
		h:mesh = "fvcom_mesh" ;
		h:location = "node" ;
	float nv(three, nele) ;
		nv:long_name = "nodes surrounding element" ;
		nv:cf_role = "face_node_connectivity" ;
		nv:start_index = 1 ;
	float zeta(time, node) ;
		zeta:long_name = "Water Surface Elevation" ;
		zeta:units = "meters" ;
		zeta:standard_name = "sea_surface_height_above_geoid" ;
		zeta:coordinates = "time lat lon" ;
		zeta:type = "data" ;
		zeta:missing_value = -999. ;
		zeta:field = "elev, scalar" ;
		zeta:mesh = "fvcom_mesh" ;
		zeta:location = "node" ;
	float ua(time, nele) ;
		ua:long_name = "Vertically Averaged x-velocity" ;
		ua:units = "meters s-1" ;
		ua:type = "data" ;
		ua:missing_value = -999. ;
		ua:field = "ua, scalar" ;
		ua:standard_name = "barotropic_eastward_sea_water_velocity" ;
		ua:coordinates = "time latc lonc" ;
		ua:mesh = "fvcom_mesh" ;
		ua:location = "face" ;
	float va(time, nele) ;
		va:long_name = "Vertically Averaged y-velocity" ;
		va:units = "meters s-1" ;
		va:type = "data" ;
		va:missing_value = -999. ;
		va:field = "va, scalar" ;
		va:standard_name = "barotropic_northward_sea_water_velocity" ;
		va:coordinates = "time latc lonc" ;
		va:mesh = "fvcom_mesh" ;
		va:location = "face" ;
	float maxele(node) ;
		maxele:long_name = "maximum water surface elevation above geoid" ;
		maxele:units = "meters" ;
		maxele:standard_name = "maximum water surface elevation" ;
		maxele:coordinates = "lat lon" ;
		maxele:valid_min = 0.276019977037 ;
		maxele:valid_max = 6.0717921 ;
		maxele:missing_value = -999. ;
		maxele:field = "elev, scalar" ;
		maxele:mesh = "fvcom_mesh" ;
		maxele:location = "node" ;
	int fvcom_mesh ;
		fvcom_mesh:cf_role = "mesh_topology" ;
		fvcom_mesh:topology_dimension = 2 ;
		fvcom_mesh:node_coordinates = "lon lat" ;
		fvcom_mesh:face_coordinates = "lonc latc" ;
		fvcom_mesh:face_node_connectivity = "nv" ;

// global attributes:
		:model = "FVCOM" ;
		:institution = "University of North Carolina" ;
		:institution = "University of Notre Dame" ;
		:Conventions = "UGRID-0.9.0" ;
		:cdm_data_type = "ugrid" ;
		:DODS.strlen = 26 ;
		:DODS.dimName = "DateStrLen" ;
		:DODS_EXTRA.Unlimited_Dimension = "time" ;
}

